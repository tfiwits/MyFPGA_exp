library ieee;
use ieee.std_logic_1164.all;

entity nul_l is
port(
		as:out std_logic
);
end nul_l;

architecture as_null of nul_l is 
begin

end as_null; 